// The use of this code requires a license file. If you lack the license file, you are prohibited to use it!

////////////////////////////////////////////////////////////////////////////////////////////////////
// Author       : Peter Cseh
// Library      : lib_cm
// Description  : Common package that defines basic data tpyes
////////////////////////////////////////////////////////////////////////////////////////////////////

`ifndef __CM_PKG_TYPE
`define __CM_PKG_TYPE

package cm_pkg_type;

    typedef byte unsigned       u8;
    typedef shortint unsigned   u16;
    typedef int unsigned        u32;
    typedef longint unsigned    u64;

endpackage

`endif