// The use of this code requires a license file. If you lack the license file, you are prohibited to use it!

////////////////////////////////////////////////////////////////////////////////////////////////////
// Author       : Peter Cseh
// Library      : Data Stream
// Description  :
////////////////////////////////////////////////////////////////////////////////////////////////////

module fifo #(
    parameter int WIDTH = 8,
    parameter int DEPTH = 8
)(
    input logic i_clk,
    input logic i_rst,


);

endmodule