// The use of this code requires a license file. If you lack the license file, you are prohibited to use it!

////////////////////////////////////////////////////////////////////////////////////////////////////
// Author       : Peter Cseh
// Library      :
// Description  :
////////////////////////////////////////////////////////////////////////////////////////////////////

import sys_pkg_type::*;
import cm_pkg::*;

module sim_cm_sort ();

////////////////////////////////////////////////////////////////////////////////////////////////////
// Initialize (Clock & Reset)
////////////////////////////////////////////////////////////////////////////////////////////////////

    // Clock
    logic clk = 1'b0;
    always #5 clk = ~clk;

    // Reset
    logic rst = 1'b0;

    task rst_dut;
        begin
            rst <= 1'b1;
            repeat(2) @ (posedge clk);
            rst <= 1'b0;
            repeat(2) @ (posedge clk);
        end
    endtask

    initial begin
        rst_dut();
    end

////////////////////////////////////////////////////////////////////////////////////////////////////
//
////////////////////////////////////////////////////////////////////////////////////////////////////

    localparam DCNT = 8;
    localparam DWIDTH = 8;

////////////////////////////////////////////////////////////////////////////////////////////////////
//
////////////////////////////////////////////////////////////////////////////////////////////////////

    logic i_vld;
    logic [DCNT - 1 : 0][DWIDTH - 1 : 0] i_data;
    logic o_vld;
    logic [DCNT - 1 : 0][DWIDTH - 1 : 0] o_data;

////////////////////////////////////////////////////////////////////////////////////////////////////
// DUT
////////////////////////////////////////////////////////////////////////////////////////////////////

    cm_sort #(
        .DCNT(DCNT),
        .DWIDTH(DWIDTH),
        .REG_CNT(1)
    ) sort (
        .i_clk(clk),
        .i_rst(rst),
        .i_vld(i_vld),
        .i_data(i_data),
        .o_vld(o_vld),
        .o_data(o_data)
    );


    // Drive
    initial begin
        i_vld = 1'b1;
        i_data = {  8'h01, 8'h03, 8'h02, 8'h05,
                    8'h00, 8'hA0, 8'h03, 8'h01};
    end


endmodule
